library IEEE;
use IEEE.std_logic_1164.ALL;
use IEEE.numeric_std.ALL;

entity logic is
	port (
		-- TODO Implement interface definition
	);
end entity logic;

architecture behav of logic is

begin
	
	-- TODO Implement logic circuit

end behav;

