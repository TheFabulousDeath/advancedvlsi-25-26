library IEEE;
use IEEE.std_logic_1164.ALL;
use IEEE.numeric_std.ALL;

entity program_counter_tb is
	generic (
		
	);
	port (
		
	);
end entity program_counter_tb;

